// -------------------- INSTRUCTION DECODER --------------------
// idk mb i aint good at this, need mo booze

`timescale 1ns/1ns

module instruction_decoder(
	input [INSTR_WIDTH-1:0] INSTRUCTION,
	output reg RESET_INSTR,
	output reg MEM_SEL,
	output reg [1:0] MUX_SEL,
	output reg CE_R0,
	output reg CE_ACC,
	output reg REG_WR,
	output reg CE_RAM,
	output reg [1:0] JUMP,
	output reg [OP_WIDTH-1:0] OP,
	output reg CE_STACK,
	output reg nRW_STACK,
	output reg STACK_SEL,
	output reg PC_SEL,
	output reg CE_PORTA
);

parameter INSTR_WIDTH = 5;
parameter OP_WIDTH = 4;

always @(*) begin
	case(INSTRUCTION)
		5'h00: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000000000101010000; // NOP
		5'h01: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000000000000010010; // NOT
		5'h02: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000000000100010010; // DEC
		5'h03: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000000000100110010; // INC
		5'h04: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000000000001010010; // OR
		5'h05: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000000000001110010; // AND
		5'h06: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000000000110010010; // XOR
		5'h07: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000000000101000000; // XNOR
		5'h08: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000000000011110010; // RL
		5'h09: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000000000011010010; // RR
		5'h0A: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000000000010110010; // ADD
		5'h0B: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000000000010010010; // SUB
		5'h0C: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000000000101000000; // ADDC (N/A)
		5'h0D: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000000000101000000; // SUBC (N/A)
		5'h0E: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000000000101000000; // LDIL (N/A)
		5'h0F: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000000000101010110; // LDI, LDIH (N/A)
		5'h10: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000000000101110010; // LD R
		5'h11: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000000000101010001; // ST R
		5'h12: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000000001101110010; // MOV A,@R
		5'h13: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000000010101010000; // MOV @R,A
		5'h14: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000110000101010000; // PUSH
		5'h15: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000100000101011010; // POP
		5'h16: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000000000101011110; // READ
		5'h17: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b100000000101010000; // WRITE
		5'h18: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b001111100101010000; // CALL
		5'h19: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b010101100101010000; // RET
		5'h1A: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000001100101010000; // JMP
		5'h1B: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000000100101010000; // JZ
		5'h1C: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000001000101010000; // JNZ
		5'h1D: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000000000101000000;
		5'h1E: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000000000101000000;
		5'h1F: {CE_PORTA, PC_SEL, STACK_SEL, CE_STACK, nRW_STACK, JUMP[1:0], CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL[1:0], CE_ACC, REG_WR} <= 18'b000000000101000000; // RST
	endcase
end

endmodule // instruction_decoder