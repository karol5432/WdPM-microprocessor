// -------------------- INSTRUCTION DECODER --------------------
// idk mb i aint good at this, need mo booze

module instruction_decoder(
	input [INSTR_WIDTH-1:0] INSTRUCTION,
	output reg RESET_INSTR,
	output reg MEM_SEL,
	output reg MUX_SEL,
	output reg CE_R0,
	output reg CE_ACC,
	output reg REG_WR,
	output reg CE_RAM,
	output reg CE_PC,
	output reg [OP_WIDTH-1:0] OP
);

parameter INSTR_WIDTH = 5;
parameter OP_WIDTH = 4;

always @(*) begin
	case(INSTRUCTION)
	//					RESET SEL CE(reg) CE(acc) inst1 inst0
		5'h00: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00000000010; // NOT
		5'h01: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00000010010; // XOR
		5'h02: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00000100010; // OR
		5'h03: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00000110010; // AND
		5'h04: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00001000010; // SUB
		5'h05: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00001010010; // ADD R
		5'h06: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00001100010; // RR
		5'h07: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00001110010; // RL
		5'h08: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00010000010; // DEC
		5'h09: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00010010010; // INC
		5'h0A: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00010110010; // LD R
		5'h0B: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00010100001; // ST R
		5'h0C: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00010100000; // NOP
		5'h0D: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00010100110; // LDI
		5'h0E: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00010101000; // RST
		5'h0F: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00010101000; // RST
		5'h10: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00110110010; // MOV A,#addr // nie zadziala, bo potrzeba 2 taktow zegarowych, mozna zrobic MOV A,@R0, ale najpierw trzeba naprawic R0 bo nie dziala
		5'h11: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b01010100000; // MOV #addr,A // nie dziala bo chyba jak sie ustawia wartosci to tylko w nastepnym takcie dzialaja, nie fajnie
		5'h12: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00000100010; // PUSH
		5'h13: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00000110010; // POP
		5'h14: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b10010100000; // JMP IMM
		5'h15: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00001010010;
		5'h16: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00001100010;
		5'h17: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00001110010;
		5'h18: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00010000010;
		5'h19: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00010010010;
		5'h1A: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00010110010;
		5'h1B: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00010100001;
		5'h1C: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00010100000;
		5'h1D: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00010100110;
		5'h1E: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00010101000;
		5'h1F: {CE_PC, CE_RAM, MEM_SEL, OP[OP_WIDTH-1:0], RESET_INSTR, MUX_SEL, CE_ACC, REG_WR} <= 11'b00010101000; // RST
	endcase
end

endmodule // instruction_decoder